module memory
    #(parameter data_width = 256,
      parameter addr_width = 16)
     (input  [addr_width-1:0] address,
      input  [data_width-1:0] data_write,
      input                   clk,
      input                   we,
      input                   reset,
      input                   petition,
      output reg              serviceReady,
      //output reg [data_width-1:0] data_read_high,
      output reg [data_width-1:0] data_read);
//we are not yet implementing the writes

    reg [data_width-1:0] mem [0:(2**addr_width)-1];
    reg [1:0] state;
    reg enable_output_register;
    wire [addr_width-1:0] previousAddress;
/*    always @(posedge clk) begin : write_proc
        if (we == 1)begin
            mem[address] = data_write_high;
            mem[address+1] = data_write_low;
        end
    end
*/

  register #(256) output_register(
    .clk(clk),
    .enable(enable_output_register), //the enable is generated by the decode itself
    .reset(reset),
    .d({mem[address+14], mem[address+12], mem[address+10], mem[address+8], mem[address+6], mem[address+4], mem[address+2], mem[address]}),
    
    .q(data_read)
  );

  register #(addr_width) address_register(
    .clk(clk),
    .enable(enable_output_register), //the enable is generated by the decode itself
    .reset(reset),
    .d(address),
    
    .q(previousAddress)
  );

    parameter zero=0, one=1, two=2, three=3;

//se necesita implementar un registro de cambio de dirección
//nos servira para cambiar de dirección. De otra manera podemos
//dar xxxx para los ciclos cuando no se leen datos utiles.
  always @(state) 
    begin
    case (state)
      zero:
      begin
        serviceReady <= 1'b0;
        enable_output_register <= 1'b0;
      end
      one:
      begin
        serviceReady <= 1'b0;
        enable_output_register <= 1'b0;
      end
      two:
      begin
        serviceReady <= 1'b0;
        enable_output_register <= 1'b1;
      end
      three:
      begin
        serviceReady <= 1'b1;
        enable_output_register <= 1'b0;
        //next cycle the instruction may advance 
        //to cache stage and have read the valid data
        //in case of instructions, serviceReady
        //cycle is needed
      end
      default:
        begin
        serviceReady = 1'b0;
        enable_output_register <= 1'b0;
        end
    endcase
  end

  always @(posedge clk or posedge reset or address)
    begin
      if (reset)
        state = zero;
      else
        if (petition)
          case (state) //petition is set to 1 in case of miss
            zero:
              if (address != previousAddress) 
                state = zero;
              else
                state = one;
            one:
              if (address != previousAddress) 
                state = zero;
              else
                state = two;
            two:
              if (address != previousAddress) 
                state = zero;
              else
                state = three;
            three:
              state = zero;
               //in the third cycle no cancelling
               //should be requested
          endcase
        else
          state = zero;
      end
endmodule
