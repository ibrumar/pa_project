module instr_cache
     #(parameter cache_line_width = 256,
      parameter word_width = 16,
      //in the data cache we will access not only
      //data with width 'word_width'
      parameter addr_width = 16,
      parameter num_cache_lines = 4)
     (
      //inputs from processor

      input  [addr_width-1:0] address,
      input                   clk,
      //inputs from arbiter
      input                   pet,
      //input from memory
      input                   dataReadFromMem,
      input                   memServiceReady,
      output
      //output to processor
      output [word_width-1:0] instructionBits,
      output                  isHit,
      //output to arbitrer
      output [addr_width-1:0] addrToArb, //we keep this
                                         //to be consistent
                                         //with the data cache
      output                  petitionToArb,
      );


//you need 4 registers x 256bits for the lines
//4 registers x 16 bits for tags -> maybe less. Compute
//how many
//you need a multiplexer for the line of 4 lines x 256 bits, and
//another multiplexer for the word of 16 words x 16 bits
//a validity bit vector is necessary. One bit per line.

   //Tags
   
   //Validity bits
   //if we had a miss, the memory service is ready, the matching cache
   //line is written
   wire                              canWriteValidity = !isHit && memServiceReady;
   wire signed [num_cache_lines-1:0] validityExtended = canWriteValidity;
   wire [num_cache_lines-1:0]        enableValidityBits = validityExtended&decodedLine;
   wire [num_cache_lines-1:0]        validityBits; //this is the output of the
   //validity register

   //DATA
      //this wires come from the data lines (registers of 256 bits)
   wire [cache_line_width-1:0] dataLines [0:num_cache_lines-1];

   reg [word_width-1:0] selectedLine [16*word_width] = dataLines[address[5:4]];
   reg [word_width-1:0] selectedWord = selectedLine[address[3:0]];
                                    
  assign addrToArb = address;
  
  reg [num_cache_lines-1:0] decodedLine;

  always @(*)
    begin
      case (address[5:4]) //those bits are the cache line
      2'b00:
        decodedLine <= 4'b0001;

      2'b01:
        decodedLine <= 4'b0010;

      2'b10:
        decodedLine <= 4'b0100;
      
      2'b11:
        decodedLine <= 4'b1000;
      endcase
    end

  genvar i;
  generate
    for (i=0; i<num_cache_lines; i=i+1)
      begin: gen_register
        register #(cache_line_width) my_register(.clk(clk),
                           .enable(decoded_line), //BAD_DONE. You enable only when the line comes from memory 
                           .reset(reset),
                           .d(dataReadFromMem)
                           .q(dataLines[i]);
      end
  endgenerate

  //validity register is set on first retrieval
  //upon on an invalid line
  register #(num_cache_lines) validity_register(
    .clk(clk),
    .enable(enable_validity_register), //the enable is generated by the decode itself
    .reset(reset),
    .d(1'b1), //you must create this reg variable
    
    .q(validityBits)
  );
 
 //for tommorrow generate the cables for the tags registers
 //and add the logic for miss. You need to modify the register enbable to
 //be active only when data comes from memory. The validity bit enable
 //is very close to this.

endmodule
